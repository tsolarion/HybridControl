-- megafunction wizard: %ALTFP_CONVERT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTFP_CONVERT 

-- ============================================================
-- File Name: fp32_signed16_conv.vhd
-- Megafunction Name(s):
-- 			ALTFP_CONVERT
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 16.1.0 Build 196 10/24/2016 SJ Standard Edition
-- ************************************************************


--Copyright (C) 2016  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel MegaCore Function License Agreement, or other 
--applicable license agreement, including, without limitation, 
--that your use is for the sole purpose of programming logic 
--devices manufactured by Intel and sold by Intel or its 
--authorized distributors.  Please refer to the applicable 
--agreement for further details.


--altfp_convert CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" OPERATION="FLOAT2FIXED" ROUNDING="TO_NEAREST" WIDTH_DATA=32 WIDTH_EXP_INPUT=8 WIDTH_EXP_OUTPUT=8 WIDTH_INT=4 WIDTH_MAN_INPUT=23 WIDTH_MAN_OUTPUT=23 WIDTH_RESULT=16 clock dataa nan overflow result underflow
--VERSION_BEGIN 16.1 cbx_altbarrel_shift 2016:10:24:15:04:16:SJ cbx_altera_syncram_nd_impl 2016:10:24:15:04:16:SJ cbx_altfp_convert 2016:10:24:15:04:16:SJ cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_altsyncram 2016:10:24:15:04:16:SJ cbx_cycloneii 2016:10:24:15:04:16:SJ cbx_lpm_abs 2016:10:24:15:04:16:SJ cbx_lpm_add_sub 2016:10:24:15:04:16:SJ cbx_lpm_compare 2016:10:24:15:04:16:SJ cbx_lpm_decode 2016:10:24:15:04:16:SJ cbx_lpm_divide 2016:10:24:15:04:16:SJ cbx_lpm_mux 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ cbx_nadder 2016:10:24:15:04:16:SJ cbx_stratix 2016:10:24:15:04:16:SJ cbx_stratixii 2016:10:24:15:04:16:SJ cbx_stratixiii 2016:10:24:15:04:16:SJ cbx_stratixv 2016:10:24:15:04:16:SJ cbx_util_mgl 2016:10:24:15:04:16:SJ  VERSION_END


--altbarrel_shift CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" PIPELINE=2 SHIFTDIR="VARIABLE" SHIFTTYPE="LOGICAL" WIDTH=38 WIDTHDIST=6 aclr clk_en clock data direction distance result
--VERSION_BEGIN 16.1 cbx_altbarrel_shift 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ  VERSION_END

--synthesis_resources = reg 81 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fp32_signed16_conv_altbarrel_shift_i4h IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clk_en	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (37 DOWNTO 0);
		 direction	:	IN  STD_LOGIC := '0';
		 distance	:	IN  STD_LOGIC_VECTOR (5 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (37 DOWNTO 0)
	 ); 
 END fp32_signed16_conv_altbarrel_shift_i4h;

 ARCHITECTURE RTL OF fp32_signed16_conv_altbarrel_shift_i4h IS

	 SIGNAL	 dir_pipe	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sbit_piper1d	:	STD_LOGIC_VECTOR(37 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sbit_piper2d	:	STD_LOGIC_VECTOR(37 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sel_pipec3r1d	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sel_pipec4r1d	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sel_pipec5r1d	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range321w333w334w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range321w329w330w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range342w354w355w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range342w350w351w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range364w376w377w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range364w372w373w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range387w398w399w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range387w394w395w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range406w417w418w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range406w413w414w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range427w438w439w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range427w434w435w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range321w325w326w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range342w346w347w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range364w368w369w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range387w390w391w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range406w409w410w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range427w430w431w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range321w333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range321w329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range342w354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range342w350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range364w376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range364w372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range387w398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range387w394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range406w417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range406w413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range427w438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range427w434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_dir_w_range318w332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_dir_w_range340w353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_dir_w_range361w375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_dir_w_range385w397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_dir_w_range404w416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_dir_w_range424w437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range321w325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range342w346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range364w368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range387w390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range406w409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range427w430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range321w333w334w335w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range342w354w355w356w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range364w376w377w378w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range387w398w399w400w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range406w417w418w419w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range427w438w439w440w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w336w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w357w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w379w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w401w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w420w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w441w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  dir_w :	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  direction_w :	STD_LOGIC;
	 SIGNAL  pad_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  sbit_w :	STD_LOGIC_VECTOR (265 DOWNTO 0);
	 SIGNAL  sel_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  smux_w :	STD_LOGIC_VECTOR (227 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w328w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w331w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w349w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w352w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w371w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w374w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w393w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w396w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w412w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w415w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w433w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w436w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_dir_w_range318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_dir_w_range340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_dir_w_range361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_dir_w_range385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_dir_w_range404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_dir_w_range424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sbit_w_range359w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sbit_w_range381w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sbit_w_range403w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sbit_w_range422w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sbit_w_range316w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sbit_w_range339w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sel_w_range321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sel_w_range342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sel_w_range364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sel_w_range387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sel_w_range406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sel_w_range427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_smux_w_range380w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_smux_w_range442w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
 BEGIN

	loop0 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range321w333w334w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range321w333w(0) AND wire_altbarrel_shift2_w331w(i);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range321w329w330w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range321w329w(0) AND wire_altbarrel_shift2_w328w(i);
	END GENERATE loop1;
	loop2 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range342w354w355w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range342w354w(0) AND wire_altbarrel_shift2_w352w(i);
	END GENERATE loop2;
	loop3 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range342w350w351w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range342w350w(0) AND wire_altbarrel_shift2_w349w(i);
	END GENERATE loop3;
	loop4 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range364w376w377w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range364w376w(0) AND wire_altbarrel_shift2_w374w(i);
	END GENERATE loop4;
	loop5 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range364w372w373w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range364w372w(0) AND wire_altbarrel_shift2_w371w(i);
	END GENERATE loop5;
	loop6 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range387w398w399w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range387w398w(0) AND wire_altbarrel_shift2_w396w(i);
	END GENERATE loop6;
	loop7 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range387w394w395w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range387w394w(0) AND wire_altbarrel_shift2_w393w(i);
	END GENERATE loop7;
	loop8 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range406w417w418w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range406w417w(0) AND wire_altbarrel_shift2_w415w(i);
	END GENERATE loop8;
	loop9 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range406w413w414w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range406w413w(0) AND wire_altbarrel_shift2_w412w(i);
	END GENERATE loop9;
	loop10 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range427w438w439w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range427w438w(0) AND wire_altbarrel_shift2_w436w(i);
	END GENERATE loop10;
	loop11 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range427w434w435w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range427w434w(0) AND wire_altbarrel_shift2_w433w(i);
	END GENERATE loop11;
	loop12 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range321w325w326w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range321w325w(0) AND wire_altbarrel_shift2_w_sbit_w_range316w(i);
	END GENERATE loop12;
	loop13 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range342w346w347w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range342w346w(0) AND wire_altbarrel_shift2_w_sbit_w_range339w(i);
	END GENERATE loop13;
	loop14 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range364w368w369w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range364w368w(0) AND wire_altbarrel_shift2_w_sbit_w_range359w(i);
	END GENERATE loop14;
	loop15 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range387w390w391w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range387w390w(0) AND wire_altbarrel_shift2_w_sbit_w_range381w(i);
	END GENERATE loop15;
	loop16 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range406w409w410w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range406w409w(0) AND wire_altbarrel_shift2_w_sbit_w_range403w(i);
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range427w430w431w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range427w430w(0) AND wire_altbarrel_shift2_w_sbit_w_range422w(i);
	END GENERATE loop17;
	wire_altbarrel_shift2_w_lg_w_sel_w_range321w333w(0) <= wire_altbarrel_shift2_w_sel_w_range321w(0) AND wire_altbarrel_shift2_w_lg_w_dir_w_range318w332w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range321w329w(0) <= wire_altbarrel_shift2_w_sel_w_range321w(0) AND wire_altbarrel_shift2_w_dir_w_range318w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range342w354w(0) <= wire_altbarrel_shift2_w_sel_w_range342w(0) AND wire_altbarrel_shift2_w_lg_w_dir_w_range340w353w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range342w350w(0) <= wire_altbarrel_shift2_w_sel_w_range342w(0) AND wire_altbarrel_shift2_w_dir_w_range340w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range364w376w(0) <= wire_altbarrel_shift2_w_sel_w_range364w(0) AND wire_altbarrel_shift2_w_lg_w_dir_w_range361w375w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range364w372w(0) <= wire_altbarrel_shift2_w_sel_w_range364w(0) AND wire_altbarrel_shift2_w_dir_w_range361w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range387w398w(0) <= wire_altbarrel_shift2_w_sel_w_range387w(0) AND wire_altbarrel_shift2_w_lg_w_dir_w_range385w397w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range387w394w(0) <= wire_altbarrel_shift2_w_sel_w_range387w(0) AND wire_altbarrel_shift2_w_dir_w_range385w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range406w417w(0) <= wire_altbarrel_shift2_w_sel_w_range406w(0) AND wire_altbarrel_shift2_w_lg_w_dir_w_range404w416w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range406w413w(0) <= wire_altbarrel_shift2_w_sel_w_range406w(0) AND wire_altbarrel_shift2_w_dir_w_range404w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range427w438w(0) <= wire_altbarrel_shift2_w_sel_w_range427w(0) AND wire_altbarrel_shift2_w_lg_w_dir_w_range424w437w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range427w434w(0) <= wire_altbarrel_shift2_w_sel_w_range427w(0) AND wire_altbarrel_shift2_w_dir_w_range424w(0);
	wire_altbarrel_shift2_w_lg_w_dir_w_range318w332w(0) <= NOT wire_altbarrel_shift2_w_dir_w_range318w(0);
	wire_altbarrel_shift2_w_lg_w_dir_w_range340w353w(0) <= NOT wire_altbarrel_shift2_w_dir_w_range340w(0);
	wire_altbarrel_shift2_w_lg_w_dir_w_range361w375w(0) <= NOT wire_altbarrel_shift2_w_dir_w_range361w(0);
	wire_altbarrel_shift2_w_lg_w_dir_w_range385w397w(0) <= NOT wire_altbarrel_shift2_w_dir_w_range385w(0);
	wire_altbarrel_shift2_w_lg_w_dir_w_range404w416w(0) <= NOT wire_altbarrel_shift2_w_dir_w_range404w(0);
	wire_altbarrel_shift2_w_lg_w_dir_w_range424w437w(0) <= NOT wire_altbarrel_shift2_w_dir_w_range424w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range321w325w(0) <= NOT wire_altbarrel_shift2_w_sel_w_range321w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range342w346w(0) <= NOT wire_altbarrel_shift2_w_sel_w_range342w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range364w368w(0) <= NOT wire_altbarrel_shift2_w_sel_w_range364w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range387w390w(0) <= NOT wire_altbarrel_shift2_w_sel_w_range387w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range406w409w(0) <= NOT wire_altbarrel_shift2_w_sel_w_range406w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range427w430w(0) <= NOT wire_altbarrel_shift2_w_sel_w_range427w(0);
	loop18 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range321w333w334w335w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range321w333w334w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range321w329w330w(i);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range342w354w355w356w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range342w354w355w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range342w350w351w(i);
	END GENERATE loop19;
	loop20 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range364w376w377w378w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range364w376w377w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range364w372w373w(i);
	END GENERATE loop20;
	loop21 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range387w398w399w400w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range387w398w399w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range387w394w395w(i);
	END GENERATE loop21;
	loop22 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range406w417w418w419w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range406w417w418w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range406w413w414w(i);
	END GENERATE loop22;
	loop23 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range427w438w439w440w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range427w438w439w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range427w434w435w(i);
	END GENERATE loop23;
	loop24 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w336w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range321w333w334w335w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range321w325w326w(i);
	END GENERATE loop24;
	loop25 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w357w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range342w354w355w356w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range342w346w347w(i);
	END GENERATE loop25;
	loop26 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w379w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range364w376w377w378w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range364w368w369w(i);
	END GENERATE loop26;
	loop27 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w401w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range387w398w399w400w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range387w390w391w(i);
	END GENERATE loop27;
	loop28 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w420w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range406w417w418w419w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range406w409w410w(i);
	END GENERATE loop28;
	loop29 : FOR i IN 0 TO 37 GENERATE 
		wire_altbarrel_shift2_w441w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range427w438w439w440w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range427w430w431w(i);
	END GENERATE loop29;
	dir_w <= ( dir_pipe(1) & dir_w(4 DOWNTO 3) & dir_pipe(0) & dir_w(1 DOWNTO 0) & direction_w);
	direction_w <= direction;
	pad_w <= (OTHERS => '0');
	result <= sbit_w(265 DOWNTO 228);
	sbit_w <= ( sbit_piper2d & smux_w(189 DOWNTO 114) & sbit_piper1d & smux_w(75 DOWNTO 0) & data);
	sel_w <= ( sel_pipec5r1d & sel_pipec4r1d & sel_pipec3r1d & distance(2 DOWNTO 0));
	smux_w <= ( wire_altbarrel_shift2_w441w & wire_altbarrel_shift2_w420w & wire_altbarrel_shift2_w401w & wire_altbarrel_shift2_w379w & wire_altbarrel_shift2_w357w & wire_altbarrel_shift2_w336w);
	wire_altbarrel_shift2_w328w <= ( pad_w(0) & sbit_w(37 DOWNTO 1));
	wire_altbarrel_shift2_w331w <= ( sbit_w(36 DOWNTO 0) & pad_w(0));
	wire_altbarrel_shift2_w349w <= ( pad_w(1 DOWNTO 0) & sbit_w(75 DOWNTO 40));
	wire_altbarrel_shift2_w352w <= ( sbit_w(73 DOWNTO 38) & pad_w(1 DOWNTO 0));
	wire_altbarrel_shift2_w371w <= ( pad_w(3 DOWNTO 0) & sbit_w(113 DOWNTO 80));
	wire_altbarrel_shift2_w374w <= ( sbit_w(109 DOWNTO 76) & pad_w(3 DOWNTO 0));
	wire_altbarrel_shift2_w393w <= ( pad_w(7 DOWNTO 0) & sbit_w(151 DOWNTO 122));
	wire_altbarrel_shift2_w396w <= ( sbit_w(143 DOWNTO 114) & pad_w(7 DOWNTO 0));
	wire_altbarrel_shift2_w412w <= ( pad_w(15 DOWNTO 0) & sbit_w(189 DOWNTO 168));
	wire_altbarrel_shift2_w415w <= ( sbit_w(173 DOWNTO 152) & pad_w(15 DOWNTO 0));
	wire_altbarrel_shift2_w433w <= ( pad_w(31 DOWNTO 0) & sbit_w(227 DOWNTO 222));
	wire_altbarrel_shift2_w436w <= ( sbit_w(195 DOWNTO 190) & pad_w(31 DOWNTO 0));
	wire_altbarrel_shift2_w_dir_w_range318w(0) <= dir_w(0);
	wire_altbarrel_shift2_w_dir_w_range340w(0) <= dir_w(1);
	wire_altbarrel_shift2_w_dir_w_range361w(0) <= dir_w(2);
	wire_altbarrel_shift2_w_dir_w_range385w(0) <= dir_w(3);
	wire_altbarrel_shift2_w_dir_w_range404w(0) <= dir_w(4);
	wire_altbarrel_shift2_w_dir_w_range424w(0) <= dir_w(5);
	wire_altbarrel_shift2_w_sbit_w_range359w <= sbit_w(113 DOWNTO 76);
	wire_altbarrel_shift2_w_sbit_w_range381w <= sbit_w(151 DOWNTO 114);
	wire_altbarrel_shift2_w_sbit_w_range403w <= sbit_w(189 DOWNTO 152);
	wire_altbarrel_shift2_w_sbit_w_range422w <= sbit_w(227 DOWNTO 190);
	wire_altbarrel_shift2_w_sbit_w_range316w <= sbit_w(37 DOWNTO 0);
	wire_altbarrel_shift2_w_sbit_w_range339w <= sbit_w(75 DOWNTO 38);
	wire_altbarrel_shift2_w_sel_w_range321w(0) <= sel_w(0);
	wire_altbarrel_shift2_w_sel_w_range342w(0) <= sel_w(1);
	wire_altbarrel_shift2_w_sel_w_range364w(0) <= sel_w(2);
	wire_altbarrel_shift2_w_sel_w_range387w(0) <= sel_w(3);
	wire_altbarrel_shift2_w_sel_w_range406w(0) <= sel_w(4);
	wire_altbarrel_shift2_w_sel_w_range427w(0) <= sel_w(5);
	wire_altbarrel_shift2_w_smux_w_range380w <= smux_w(113 DOWNTO 76);
	wire_altbarrel_shift2_w_smux_w_range442w <= smux_w(227 DOWNTO 190);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dir_pipe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dir_pipe <= ( dir_w(5) & dir_w(2));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sbit_piper1d <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sbit_piper1d <= wire_altbarrel_shift2_w_smux_w_range380w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sbit_piper2d <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sbit_piper2d <= wire_altbarrel_shift2_w_smux_w_range442w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sel_pipec3r1d <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sel_pipec3r1d <= distance(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sel_pipec4r1d <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sel_pipec4r1d <= distance(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sel_pipec5r1d <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sel_pipec5r1d <= distance(5);
			END IF;
		END IF;
	END PROCESS;

 END RTL; --fp32_signed16_conv_altbarrel_shift_i4h

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 6 lpm_compare 4 reg 226 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fp32_signed16_conv_altfp_convert_46p IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 dataa	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 nan	:	OUT  STD_LOGIC;
		 overflow	:	OUT  STD_LOGIC;
		 result	:	OUT  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 underflow	:	OUT  STD_LOGIC
	 ); 
 END fp32_signed16_conv_altfp_convert_46p;

 ARCHITECTURE RTL OF fp32_signed16_conv_altfp_convert_46p IS

	 SIGNAL  wire_altbarrel_shift2_distance	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_barrel_direction_negative164w165w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_result	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL	 added_power2_reg	:	STD_LOGIC_VECTOR(5 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_direction_negative_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 below_lower_limit2_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 below_lower_limit2_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 below_lower_limit2_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 below_lower_limit2_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_below_lower_limit2_reg4_w_lg_q288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 below_lower_limit3_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 below_lower_limit3_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 below_lower_limit3_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 below_lower_limit3_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_below_lower_limit3_reg4_w_lg_q292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 border_lower_limit_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 border_lower_limit_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 border_lower_limit_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 border_lower_limit_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_border_lower_limit_reg4_w_lg_q287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dataa_reg	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 equal_upper_limit_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 equal_upper_limit_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 equal_upper_limit_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_equal_upper_limit_reg3_w_lg_q252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 exceed_upper_limit_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exceed_upper_limit_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exceed_upper_limit_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_exceed_upper_limit_reg3_w_lg_q253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 exceed_upper_limit_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_and_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_and_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_and_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_and_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_or_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_or_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_or_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_or_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_exp_or_reg4_w_lg_q118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 int_or1_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 int_or2_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 int_or_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 int_or_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_int_or_reg3_w_lg_q251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 integer_result_reg	:	STD_LOGIC_VECTOR(15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 integer_rounded_reg	:	STD_LOGIC_VECTOR(14 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lowest_int_sel_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_lowest_int_sel_reg_w_lg_q289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 man_or1_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_or2_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_or_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_or_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_or_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_man_or_reg4_w_lg_q120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 mantissa_input_reg	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 max_shift_exceeder_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 max_shift_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 overflow_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 power2_value_reg	:	STD_LOGIC_VECTOR(5 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_input_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_input_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_input_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_sign_input_reg3_w_lg_q254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_sign_input_reg3_w_lg_q256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 sign_input_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 underflow_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_add_1_adder_cout	:	STD_LOGIC;
	 SIGNAL  wire_add_1_adder_datab	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_add_1_adder_result	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_add_sub1_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_add_sub1_result	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_add_sub3_w_lg_w_lg_cout263w264w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_add_sub3_w_lg_cout262w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_add_sub3_w_lg_cout263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub3_cout	:	STD_LOGIC;
	 SIGNAL  wire_add_sub3_datab	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_add_sub3_result	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_add_sub4_datab	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_add_sub4_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_barrel_direction_invert_dataa	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_barrel_direction_invert_result	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_power2_value_w_lg_w_result_range146w154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_power2_value_w_lg_w_lg_w_result_range146w154w155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_power2_value_overflow	:	STD_LOGIC;
	 SIGNAL  wire_power2_value_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_power2_value_w_result_range128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_power2_value_w_result_range131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_power2_value_w_result_range134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_power2_value_w_result_range137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_power2_value_w_result_range140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_power2_value_w_result_range143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_power2_value_w_result_range146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_below_lower_limit1_aeb	:	STD_LOGIC;
	 SIGNAL  wire_below_lower_limit2_aeb	:	STD_LOGIC;
	 SIGNAL  wire_below_lower_limit2_alb	:	STD_LOGIC;
	 SIGNAL  wire_exceed_upper_limit_aeb	:	STD_LOGIC;
	 SIGNAL  wire_exceed_upper_limit_agb	:	STD_LOGIC;
	 SIGNAL  wire_max_shift_compare_agb	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_add_1_w239w240w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_barrel_direction_negative162w163w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_below_limit_exceeders301w302w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_exceed_limit_exceeders312w313w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_lowest_integer_selector245w246w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_sign_input_w268w305w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_sign_input_w268w269w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_w_lg_add_1_w238w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_w_lg_barrel_direction_negative164w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_w_lg_below_limit_exceeders300w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_exceed_limit_exceeders311w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_lowest_integer_selector244w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_w_lg_sign_input_w304w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_sign_input_w267w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_below_lower_limit3_anding_range126w129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_below_lower_limit3_anding_range130w132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_below_lower_limit3_anding_range133w135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_below_lower_limit3_anding_range136w138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_below_lower_limit3_anding_range139w141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_below_lower_limit3_anding_range142w144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_below_lower_limit3_anding_range145w147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range8w13w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range14w18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range19w23w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range24w28w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range29w33w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range34w38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range39w43w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_add_1_w239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_barrel_direction_negative162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_below_limit_exceeders301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_denormal_input_w290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exceed_limit_exceeders312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_lowest_integer_selector245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_nan_input_w307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sign_input_w268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_zero_input_w291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_denormal_input_w296w297w298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_denormal_input_w296w297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_infinity_input_w308w309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_denormal_input_w296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_infinity_input_w308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_below_lower_limit3_oring_range149w151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range6w11w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range12w16w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range17w21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range22w26w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range27w31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range32w36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range37w41w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range47w50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range75w77w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range72w74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range69w71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range66w68w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range63w65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range60w62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range57w59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range54w56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range51w53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range85w87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range81w84w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range112w114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range109w111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range106w108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range103w105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range100w102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range97w99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range94w96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range91w93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range88w90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range171w174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range202w204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range205w207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range208w210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range211w213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range214w216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range217w219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range220w222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range223w225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range226w228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range229w231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range175w177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range232w234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range178w180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range181w183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range184w186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range187w189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range190w192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range193w195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range196w198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range199w201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  aclr	:	STD_LOGIC;
	 SIGNAL  add_1_cout_w :	STD_LOGIC;
	 SIGNAL  add_1_w :	STD_LOGIC;
	 SIGNAL  all_zeroes_w :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  barrel_direction_negative :	STD_LOGIC;
	 SIGNAL  barrel_mantissa_input :	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  barrel_zero_padding_w :	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  below_limit_exceeders :	STD_LOGIC;
	 SIGNAL  below_limit_integer :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  below_lower_limit2_w :	STD_LOGIC;
	 SIGNAL  below_lower_limit3_anding :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  below_lower_limit3_oring :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  below_lower_limit3_w :	STD_LOGIC;
	 SIGNAL  bias_value_less_1_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  const_bias_value_add_width_res_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  denormal_input_w :	STD_LOGIC;
	 SIGNAL  equal_upper_limit_w :	STD_LOGIC;
	 SIGNAL  exceed_limit_exceeders :	STD_LOGIC;
	 SIGNAL  exceed_limit_integer :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  exceed_upper_limit_w :	STD_LOGIC;
	 SIGNAL  exp_and :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_and_w :	STD_LOGIC;
	 SIGNAL  exp_bus :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_or :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_or_w :	STD_LOGIC;
	 SIGNAL  exponent_input :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  guard_bit_w :	STD_LOGIC;
	 SIGNAL  implied_mantissa_input :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  infinity_input_w :	STD_LOGIC;
	 SIGNAL  infinity_value_w :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  int_or1_w :	STD_LOGIC;
	 SIGNAL  int_or2_w :	STD_LOGIC;
	 SIGNAL  integer_output :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  integer_post_round :	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  integer_pre_round :	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  integer_result :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  integer_rounded :	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  integer_rounded_tmp :	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  integer_tmp_output :	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  inv_add_1_adder1_w :	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  inv_add_1_adder2_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  inv_integer :	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  lbarrel_shift_result_w :	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  lbarrel_shift_w :	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  lower_limit_selector :	STD_LOGIC;
	 SIGNAL  lowest_integer_selector :	STD_LOGIC;
	 SIGNAL  lowest_integer_value :	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  man_bus1 :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  man_bus2 :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  man_or1 :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  man_or1_w :	STD_LOGIC;
	 SIGNAL  man_or2 :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  man_or2_w :	STD_LOGIC;
	 SIGNAL  man_or_w :	STD_LOGIC;
	 SIGNAL  mantissa_input :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  max_shift_reg_w :	STD_LOGIC;
	 SIGNAL  max_shift_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  more_than_max_shift_w :	STD_LOGIC;
	 SIGNAL  nan_input_w :	STD_LOGIC;
	 SIGNAL  neg_infi_w :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  padded_exponent_input :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  pos_infi_w :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  power2_value_overflow_w :	STD_LOGIC;
	 SIGNAL  power2_value_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  round_bit_w :	STD_LOGIC;
	 SIGNAL  shift_value_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  sign_input :	STD_LOGIC;
	 SIGNAL  sign_input_w :	STD_LOGIC;
	 SIGNAL  signed_integer :	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  sticky_bit_w :	STD_LOGIC;
	 SIGNAL  sticky_bus :	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  sticky_or :	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  unsigned_integer :	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  upper_limit_w :	STD_LOGIC;
	 SIGNAL  zero_input_w :	STD_LOGIC;
	 SIGNAL  wire_w_below_lower_limit3_anding_range126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_below_lower_limit3_anding_range130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_below_lower_limit3_anding_range133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_below_lower_limit3_anding_range136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_below_lower_limit3_anding_range139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_below_lower_limit3_anding_range142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_below_lower_limit3_anding_range145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_below_lower_limit3_oring_range149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_below_lower_limit3_oring_range152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range8w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range14w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range19w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range24w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range29w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range34w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range10w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range15w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range20w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range25w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range30w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range35w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range6w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range12w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range22w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range27w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range32w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range37w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_inv_integer_range250w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range76w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range73w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range64w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range83w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range95w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range92w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range86w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range75w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range72w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range66w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range81w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range88w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  fp32_signed16_conv_altbarrel_shift_i4h
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clk_en	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(37 DOWNTO 0);
		direction	:	IN  STD_LOGIC := '0';
		distance	:	IN  STD_LOGIC_VECTOR(5 DOWNTO 0);
		result	:	OUT  STD_LOGIC_VECTOR(37 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	loop30 : FOR i IN 0 TO 14 GENERATE 
		wire_w_lg_w_lg_add_1_w239w240w(i) <= wire_w_lg_add_1_w239w(0) AND integer_pre_round(i);
	END GENERATE loop30;
	loop31 : FOR i IN 0 TO 5 GENERATE 
		wire_w_lg_w_lg_barrel_direction_negative162w163w(i) <= wire_w_lg_barrel_direction_negative162w(0) AND power2_value_reg(i);
	END GENERATE loop31;
	loop32 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_below_limit_exceeders301w302w(i) <= wire_w_lg_below_limit_exceeders301w(0) AND integer_output(i);
	END GENERATE loop32;
	loop33 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_exceed_limit_exceeders312w313w(i) <= wire_w_lg_exceed_limit_exceeders312w(0) AND below_limit_integer(i);
	END GENERATE loop33;
	loop34 : FOR i IN 0 TO 14 GENERATE 
		wire_w_lg_w_lg_lowest_integer_selector245w246w(i) <= wire_w_lg_lowest_integer_selector245w(0) AND integer_rounded_tmp(i);
	END GENERATE loop34;
	loop35 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_sign_input_w268w305w(i) <= wire_w_lg_sign_input_w268w(0) AND pos_infi_w(i);
	END GENERATE loop35;
	loop36 : FOR i IN 0 TO 14 GENERATE 
		wire_w_lg_w_lg_sign_input_w268w269w(i) <= wire_w_lg_sign_input_w268w(0) AND unsigned_integer(i);
	END GENERATE loop36;
	loop37 : FOR i IN 0 TO 14 GENERATE 
		wire_w_lg_add_1_w238w(i) <= add_1_w AND integer_post_round(i);
	END GENERATE loop37;
	loop38 : FOR i IN 0 TO 5 GENERATE 
		wire_w_lg_barrel_direction_negative164w(i) <= barrel_direction_negative AND wire_barrel_direction_invert_result(i);
	END GENERATE loop38;
	loop39 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_below_limit_exceeders300w(i) <= below_limit_exceeders AND all_zeroes_w(i);
	END GENERATE loop39;
	loop40 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_exceed_limit_exceeders311w(i) <= exceed_limit_exceeders AND infinity_value_w(i);
	END GENERATE loop40;
	loop41 : FOR i IN 0 TO 14 GENERATE 
		wire_w_lg_lowest_integer_selector244w(i) <= lowest_integer_selector AND lowest_integer_value(i);
	END GENERATE loop41;
	loop42 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_sign_input_w304w(i) <= sign_input_w AND neg_infi_w(i);
	END GENERATE loop42;
	loop43 : FOR i IN 0 TO 14 GENERATE 
		wire_w_lg_sign_input_w267w(i) <= sign_input_w AND signed_integer(i);
	END GENERATE loop43;
	wire_w_lg_w_below_lower_limit3_anding_range126w129w(0) <= wire_w_below_lower_limit3_anding_range126w(0) AND wire_power2_value_w_result_range128w(0);
	wire_w_lg_w_below_lower_limit3_anding_range130w132w(0) <= wire_w_below_lower_limit3_anding_range130w(0) AND wire_power2_value_w_result_range131w(0);
	wire_w_lg_w_below_lower_limit3_anding_range133w135w(0) <= wire_w_below_lower_limit3_anding_range133w(0) AND wire_power2_value_w_result_range134w(0);
	wire_w_lg_w_below_lower_limit3_anding_range136w138w(0) <= wire_w_below_lower_limit3_anding_range136w(0) AND wire_power2_value_w_result_range137w(0);
	wire_w_lg_w_below_lower_limit3_anding_range139w141w(0) <= wire_w_below_lower_limit3_anding_range139w(0) AND wire_power2_value_w_result_range140w(0);
	wire_w_lg_w_below_lower_limit3_anding_range142w144w(0) <= wire_w_below_lower_limit3_anding_range142w(0) AND wire_power2_value_w_result_range143w(0);
	wire_w_lg_w_below_lower_limit3_anding_range145w147w(0) <= wire_w_below_lower_limit3_anding_range145w(0) AND wire_power2_value_w_result_range146w(0);
	wire_w_lg_w_exp_and_range8w13w(0) <= wire_w_exp_and_range8w(0) AND wire_w_exp_bus_range10w(0);
	wire_w_lg_w_exp_and_range14w18w(0) <= wire_w_exp_and_range14w(0) AND wire_w_exp_bus_range15w(0);
	wire_w_lg_w_exp_and_range19w23w(0) <= wire_w_exp_and_range19w(0) AND wire_w_exp_bus_range20w(0);
	wire_w_lg_w_exp_and_range24w28w(0) <= wire_w_exp_and_range24w(0) AND wire_w_exp_bus_range25w(0);
	wire_w_lg_w_exp_and_range29w33w(0) <= wire_w_exp_and_range29w(0) AND wire_w_exp_bus_range30w(0);
	wire_w_lg_w_exp_and_range34w38w(0) <= wire_w_exp_and_range34w(0) AND wire_w_exp_bus_range35w(0);
	wire_w_lg_w_exp_and_range39w43w(0) <= wire_w_exp_and_range39w(0) AND wire_w_exp_bus_range40w(0);
	wire_w_lg_add_1_w239w(0) <= NOT add_1_w;
	wire_w_lg_barrel_direction_negative162w(0) <= NOT barrel_direction_negative;
	wire_w_lg_below_limit_exceeders301w(0) <= NOT below_limit_exceeders;
	wire_w_lg_denormal_input_w290w(0) <= NOT denormal_input_w;
	wire_w_lg_exceed_limit_exceeders312w(0) <= NOT exceed_limit_exceeders;
	wire_w_lg_lowest_integer_selector245w(0) <= NOT lowest_integer_selector;
	wire_w_lg_nan_input_w307w(0) <= NOT nan_input_w;
	wire_w_lg_sign_input_w268w(0) <= NOT sign_input_w;
	wire_w_lg_zero_input_w291w(0) <= NOT zero_input_w;
	wire_w_lg_w_lg_w_lg_denormal_input_w296w297w298w(0) <= wire_w_lg_w_lg_denormal_input_w296w297w(0) OR below_lower_limit3_reg4;
	wire_w_lg_w_lg_denormal_input_w296w297w(0) <= wire_w_lg_denormal_input_w296w(0) OR nan_input_w;
	wire_w_lg_w_lg_infinity_input_w308w309w(0) <= wire_w_lg_infinity_input_w308w(0) OR exceed_upper_limit_reg4;
	wire_w_lg_denormal_input_w296w(0) <= denormal_input_w OR zero_input_w;
	wire_w_lg_infinity_input_w308w(0) <= infinity_input_w OR max_shift_exceeder_reg;
	wire_w_lg_w_below_lower_limit3_oring_range149w151w(0) <= wire_w_below_lower_limit3_oring_range149w(0) OR wire_power2_value_w_result_range146w(0);
	wire_w_lg_w_exp_or_range6w11w(0) <= wire_w_exp_or_range6w(0) OR wire_w_exp_bus_range10w(0);
	wire_w_lg_w_exp_or_range12w16w(0) <= wire_w_exp_or_range12w(0) OR wire_w_exp_bus_range15w(0);
	wire_w_lg_w_exp_or_range17w21w(0) <= wire_w_exp_or_range17w(0) OR wire_w_exp_bus_range20w(0);
	wire_w_lg_w_exp_or_range22w26w(0) <= wire_w_exp_or_range22w(0) OR wire_w_exp_bus_range25w(0);
	wire_w_lg_w_exp_or_range27w31w(0) <= wire_w_exp_or_range27w(0) OR wire_w_exp_bus_range30w(0);
	wire_w_lg_w_exp_or_range32w36w(0) <= wire_w_exp_or_range32w(0) OR wire_w_exp_bus_range35w(0);
	wire_w_lg_w_exp_or_range37w41w(0) <= wire_w_exp_or_range37w(0) OR wire_w_exp_bus_range40w(0);
	wire_w_lg_w_man_or1_range47w50w(0) <= wire_w_man_or1_range47w(0) OR wire_w_man_bus1_range49w(0);
	wire_w_lg_w_man_or1_range75w77w(0) <= wire_w_man_or1_range75w(0) OR wire_w_man_bus1_range76w(0);
	wire_w_lg_w_man_or1_range72w74w(0) <= wire_w_man_or1_range72w(0) OR wire_w_man_bus1_range73w(0);
	wire_w_lg_w_man_or1_range69w71w(0) <= wire_w_man_or1_range69w(0) OR wire_w_man_bus1_range70w(0);
	wire_w_lg_w_man_or1_range66w68w(0) <= wire_w_man_or1_range66w(0) OR wire_w_man_bus1_range67w(0);
	wire_w_lg_w_man_or1_range63w65w(0) <= wire_w_man_or1_range63w(0) OR wire_w_man_bus1_range64w(0);
	wire_w_lg_w_man_or1_range60w62w(0) <= wire_w_man_or1_range60w(0) OR wire_w_man_bus1_range61w(0);
	wire_w_lg_w_man_or1_range57w59w(0) <= wire_w_man_or1_range57w(0) OR wire_w_man_bus1_range58w(0);
	wire_w_lg_w_man_or1_range54w56w(0) <= wire_w_man_or1_range54w(0) OR wire_w_man_bus1_range55w(0);
	wire_w_lg_w_man_or1_range51w53w(0) <= wire_w_man_or1_range51w(0) OR wire_w_man_bus1_range52w(0);
	wire_w_lg_w_man_or2_range85w87w(0) <= wire_w_man_or2_range85w(0) OR wire_w_man_bus2_range86w(0);
	wire_w_lg_w_man_or2_range81w84w(0) <= wire_w_man_or2_range81w(0) OR wire_w_man_bus2_range83w(0);
	wire_w_lg_w_man_or2_range112w114w(0) <= wire_w_man_or2_range112w(0) OR wire_w_man_bus2_range113w(0);
	wire_w_lg_w_man_or2_range109w111w(0) <= wire_w_man_or2_range109w(0) OR wire_w_man_bus2_range110w(0);
	wire_w_lg_w_man_or2_range106w108w(0) <= wire_w_man_or2_range106w(0) OR wire_w_man_bus2_range107w(0);
	wire_w_lg_w_man_or2_range103w105w(0) <= wire_w_man_or2_range103w(0) OR wire_w_man_bus2_range104w(0);
	wire_w_lg_w_man_or2_range100w102w(0) <= wire_w_man_or2_range100w(0) OR wire_w_man_bus2_range101w(0);
	wire_w_lg_w_man_or2_range97w99w(0) <= wire_w_man_or2_range97w(0) OR wire_w_man_bus2_range98w(0);
	wire_w_lg_w_man_or2_range94w96w(0) <= wire_w_man_or2_range94w(0) OR wire_w_man_bus2_range95w(0);
	wire_w_lg_w_man_or2_range91w93w(0) <= wire_w_man_or2_range91w(0) OR wire_w_man_bus2_range92w(0);
	wire_w_lg_w_man_or2_range88w90w(0) <= wire_w_man_or2_range88w(0) OR wire_w_man_bus2_range89w(0);
	wire_w_lg_w_sticky_or_range171w174w(0) <= wire_w_sticky_or_range171w(0) OR wire_w_sticky_bus_range173w(0);
	wire_w_lg_w_sticky_or_range202w204w(0) <= wire_w_sticky_or_range202w(0) OR wire_w_sticky_bus_range203w(0);
	wire_w_lg_w_sticky_or_range205w207w(0) <= wire_w_sticky_or_range205w(0) OR wire_w_sticky_bus_range206w(0);
	wire_w_lg_w_sticky_or_range208w210w(0) <= wire_w_sticky_or_range208w(0) OR wire_w_sticky_bus_range209w(0);
	wire_w_lg_w_sticky_or_range211w213w(0) <= wire_w_sticky_or_range211w(0) OR wire_w_sticky_bus_range212w(0);
	wire_w_lg_w_sticky_or_range214w216w(0) <= wire_w_sticky_or_range214w(0) OR wire_w_sticky_bus_range215w(0);
	wire_w_lg_w_sticky_or_range217w219w(0) <= wire_w_sticky_or_range217w(0) OR wire_w_sticky_bus_range218w(0);
	wire_w_lg_w_sticky_or_range220w222w(0) <= wire_w_sticky_or_range220w(0) OR wire_w_sticky_bus_range221w(0);
	wire_w_lg_w_sticky_or_range223w225w(0) <= wire_w_sticky_or_range223w(0) OR wire_w_sticky_bus_range224w(0);
	wire_w_lg_w_sticky_or_range226w228w(0) <= wire_w_sticky_or_range226w(0) OR wire_w_sticky_bus_range227w(0);
	wire_w_lg_w_sticky_or_range229w231w(0) <= wire_w_sticky_or_range229w(0) OR wire_w_sticky_bus_range230w(0);
	wire_w_lg_w_sticky_or_range175w177w(0) <= wire_w_sticky_or_range175w(0) OR wire_w_sticky_bus_range176w(0);
	wire_w_lg_w_sticky_or_range232w234w(0) <= wire_w_sticky_or_range232w(0) OR wire_w_sticky_bus_range233w(0);
	wire_w_lg_w_sticky_or_range178w180w(0) <= wire_w_sticky_or_range178w(0) OR wire_w_sticky_bus_range179w(0);
	wire_w_lg_w_sticky_or_range181w183w(0) <= wire_w_sticky_or_range181w(0) OR wire_w_sticky_bus_range182w(0);
	wire_w_lg_w_sticky_or_range184w186w(0) <= wire_w_sticky_or_range184w(0) OR wire_w_sticky_bus_range185w(0);
	wire_w_lg_w_sticky_or_range187w189w(0) <= wire_w_sticky_or_range187w(0) OR wire_w_sticky_bus_range188w(0);
	wire_w_lg_w_sticky_or_range190w192w(0) <= wire_w_sticky_or_range190w(0) OR wire_w_sticky_bus_range191w(0);
	wire_w_lg_w_sticky_or_range193w195w(0) <= wire_w_sticky_or_range193w(0) OR wire_w_sticky_bus_range194w(0);
	wire_w_lg_w_sticky_or_range196w198w(0) <= wire_w_sticky_or_range196w(0) OR wire_w_sticky_bus_range197w(0);
	wire_w_lg_w_sticky_or_range199w201w(0) <= wire_w_sticky_or_range199w(0) OR wire_w_sticky_bus_range200w(0);
	aclr <= '0';
	add_1_cout_w <= ((wire_add_1_adder_cout AND add_1_w) AND wire_sign_input_reg3_w_lg_q256w(0));
	add_1_w <= (round_bit_w AND (guard_bit_w OR sticky_bit_w));
	all_zeroes_w <= ( "0" & "000000000000000");
	barrel_direction_negative <= barrel_direction_negative_reg;
	barrel_mantissa_input <= ( barrel_zero_padding_w & implied_mantissa_input);
	barrel_zero_padding_w <= (OTHERS => '0');
	below_limit_exceeders <= (wire_w_lg_w_lg_w_lg_denormal_input_w296w297w298w(0) AND wire_border_lower_limit_reg4_w_lg_q287w(0));
	below_limit_integer <= (wire_w_lg_w_lg_below_limit_exceeders301w302w OR wire_w_lg_below_limit_exceeders300w);
	below_lower_limit2_w <= wire_below_lower_limit2_alb;
	below_lower_limit3_anding <= ( wire_w_lg_w_below_lower_limit3_anding_range145w147w & wire_w_lg_w_below_lower_limit3_anding_range142w144w & wire_w_lg_w_below_lower_limit3_anding_range139w141w & wire_w_lg_w_below_lower_limit3_anding_range136w138w & wire_w_lg_w_below_lower_limit3_anding_range133w135w & wire_w_lg_w_below_lower_limit3_anding_range130w132w & wire_w_lg_w_below_lower_limit3_anding_range126w129w & wire_power2_value_result(0));
	below_lower_limit3_oring <= ( wire_w_lg_w_below_lower_limit3_oring_range149w151w & wire_power2_value_result(6));
	below_lower_limit3_w <= (wire_power2_value_w_lg_w_lg_w_result_range146w154w155w(0) AND (NOT below_lower_limit3_anding(7)));
	bias_value_less_1_w <= "01111110";
	clk_en <= '1';
	const_bias_value_add_width_res_w <= "10000010";
	denormal_input_w <= (wire_exp_or_reg4_w_lg_q118w(0) AND man_or_reg4);
	equal_upper_limit_w <= wire_exceed_upper_limit_aeb;
	exceed_limit_exceeders <= (wire_w_lg_w_lg_infinity_input_w308w309w(0) AND wire_w_lg_nan_input_w307w(0));
	exceed_limit_integer <= (wire_w_lg_w_lg_exceed_limit_exceeders312w313w OR wire_w_lg_exceed_limit_exceeders311w);
	exceed_upper_limit_w <= wire_exceed_upper_limit_agb;
	exp_and <= ( wire_w_lg_w_exp_and_range39w43w & wire_w_lg_w_exp_and_range34w38w & wire_w_lg_w_exp_and_range29w33w & wire_w_lg_w_exp_and_range24w28w & wire_w_lg_w_exp_and_range19w23w & wire_w_lg_w_exp_and_range14w18w & wire_w_lg_w_exp_and_range8w13w & exp_bus(0));
	exp_and_w <= exp_and(7);
	exp_bus <= exponent_input;
	exp_or <= ( wire_w_lg_w_exp_or_range37w41w & wire_w_lg_w_exp_or_range32w36w & wire_w_lg_w_exp_or_range27w31w & wire_w_lg_w_exp_or_range22w26w & wire_w_lg_w_exp_or_range17w21w & wire_w_lg_w_exp_or_range12w16w & wire_w_lg_w_exp_or_range6w11w & exp_bus(0));
	exp_or_w <= exp_or(7);
	exponent_input <= dataa_reg(30 DOWNTO 23);
	guard_bit_w <= wire_altbarrel_shift2_result(23);
	implied_mantissa_input <= ( "1" & mantissa_input_reg);
	infinity_input_w <= (exp_and_reg4 AND wire_man_or_reg4_w_lg_q120w(0));
	infinity_value_w <= (wire_w_lg_w_lg_sign_input_w268w305w OR wire_w_lg_sign_input_w304w);
	int_or1_w <= man_or2(0);
	int_or2_w <= man_or1(8);
	integer_output <= ( sign_input_w & integer_tmp_output);
	integer_post_round <= wire_add_1_adder_result;
	integer_pre_round <= lbarrel_shift_w;
	integer_result <= exceed_limit_integer;
	integer_rounded <= (wire_w_lg_w_lg_lowest_integer_selector245w246w OR wire_w_lg_lowest_integer_selector244w);
	integer_rounded_tmp <= (wire_w_lg_w_lg_add_1_w239w240w OR wire_w_lg_add_1_w238w);
	integer_tmp_output <= (wire_w_lg_w_lg_sign_input_w268w269w OR wire_w_lg_sign_input_w267w);
	inv_add_1_adder1_w <= wire_add_sub3_result;
	inv_add_1_adder2_w <= (wire_add_sub3_w_lg_w_lg_cout263w264w OR wire_add_sub3_w_lg_cout262w);
	inv_integer <= (NOT integer_rounded_reg);
	lbarrel_shift_result_w <= wire_altbarrel_shift2_result;
	lbarrel_shift_w <= lbarrel_shift_result_w(37 DOWNTO 23);
	lower_limit_selector <= (((wire_below_lower_limit3_reg4_w_lg_q292w(0) AND wire_w_lg_denormal_input_w290w(0)) AND wire_lowest_int_sel_reg_w_lg_q289w(0)) AND wire_below_lower_limit2_reg4_w_lg_q288w(0));
	lowest_integer_selector <= '0';
	lowest_integer_value <= ( barrel_zero_padding_w & "1");
	man_bus1 <= mantissa_input(10 DOWNTO 0);
	man_bus2 <= mantissa_input(22 DOWNTO 11);
	man_or1 <= ( man_bus1(10) & wire_w_lg_w_man_or1_range47w50w & wire_w_lg_w_man_or1_range51w53w & wire_w_lg_w_man_or1_range54w56w & wire_w_lg_w_man_or1_range57w59w & wire_w_lg_w_man_or1_range60w62w & wire_w_lg_w_man_or1_range63w65w & wire_w_lg_w_man_or1_range66w68w & wire_w_lg_w_man_or1_range69w71w & wire_w_lg_w_man_or1_range72w74w & wire_w_lg_w_man_or1_range75w77w);
	man_or1_w <= man_or1(0);
	man_or2 <= ( man_bus2(11) & wire_w_lg_w_man_or2_range81w84w & wire_w_lg_w_man_or2_range85w87w & wire_w_lg_w_man_or2_range88w90w & wire_w_lg_w_man_or2_range91w93w & wire_w_lg_w_man_or2_range94w96w & wire_w_lg_w_man_or2_range97w99w & wire_w_lg_w_man_or2_range100w102w & wire_w_lg_w_man_or2_range103w105w & wire_w_lg_w_man_or2_range106w108w & wire_w_lg_w_man_or2_range109w111w & wire_w_lg_w_man_or2_range112w114w);
	man_or2_w <= man_or2(0);
	man_or_w <= (man_or1_reg1 OR man_or2_reg1);
	mantissa_input <= dataa_reg(22 DOWNTO 0);
	max_shift_reg_w <= max_shift_reg;
	max_shift_w <= "000010";
	more_than_max_shift_w <= (max_shift_reg_w AND add_1_cout_w);
	nan <= nan_reg;
	nan_input_w <= (exp_and_reg4 AND man_or_reg4);
	neg_infi_w <= ( "1" & "000000000000000");
	overflow <= overflow_reg;
	padded_exponent_input <= exponent_input;
	pos_infi_w <= ( "0" & "111111111111111");
	power2_value_overflow_w <= wire_power2_value_overflow;
	power2_value_w <= wire_power2_value_result(5 DOWNTO 0);
	result <= result_w;
	result_w <= integer_result_reg;
	round_bit_w <= wire_altbarrel_shift2_result(22);
	shift_value_w <= "01110011";
	sign_input <= dataa_reg(31);
	sign_input_w <= sign_input_reg4;
	signed_integer <= ( inv_add_1_adder2_w & inv_add_1_adder1_w);
	sticky_bit_w <= sticky_or(21);
	sticky_bus <= wire_altbarrel_shift2_result(21 DOWNTO 0);
	sticky_or <= ( wire_w_lg_w_sticky_or_range232w234w & wire_w_lg_w_sticky_or_range229w231w & wire_w_lg_w_sticky_or_range226w228w & wire_w_lg_w_sticky_or_range223w225w & wire_w_lg_w_sticky_or_range220w222w & wire_w_lg_w_sticky_or_range217w219w & wire_w_lg_w_sticky_or_range214w216w & wire_w_lg_w_sticky_or_range211w213w & wire_w_lg_w_sticky_or_range208w210w & wire_w_lg_w_sticky_or_range205w207w & wire_w_lg_w_sticky_or_range202w204w & wire_w_lg_w_sticky_or_range199w201w & wire_w_lg_w_sticky_or_range196w198w & wire_w_lg_w_sticky_or_range193w195w & wire_w_lg_w_sticky_or_range190w192w & wire_w_lg_w_sticky_or_range187w189w & wire_w_lg_w_sticky_or_range184w186w & wire_w_lg_w_sticky_or_range181w183w & wire_w_lg_w_sticky_or_range178w180w & wire_w_lg_w_sticky_or_range175w177w & wire_w_lg_w_sticky_or_range171w174w & sticky_bus(0));
	underflow <= underflow_reg;
	unsigned_integer <= integer_rounded_reg;
	upper_limit_w <= ((wire_sign_input_reg3_w_lg_q256w(0) AND (exceed_upper_limit_reg3 OR equal_upper_limit_reg3)) OR wire_sign_input_reg3_w_lg_q254w(0));
	zero_input_w <= (wire_exp_or_reg4_w_lg_q118w(0) AND wire_man_or_reg4_w_lg_q120w(0));
	wire_w_below_lower_limit3_anding_range126w(0) <= below_lower_limit3_anding(0);
	wire_w_below_lower_limit3_anding_range130w(0) <= below_lower_limit3_anding(1);
	wire_w_below_lower_limit3_anding_range133w(0) <= below_lower_limit3_anding(2);
	wire_w_below_lower_limit3_anding_range136w(0) <= below_lower_limit3_anding(3);
	wire_w_below_lower_limit3_anding_range139w(0) <= below_lower_limit3_anding(4);
	wire_w_below_lower_limit3_anding_range142w(0) <= below_lower_limit3_anding(5);
	wire_w_below_lower_limit3_anding_range145w(0) <= below_lower_limit3_anding(6);
	wire_w_below_lower_limit3_oring_range149w(0) <= below_lower_limit3_oring(0);
	wire_w_below_lower_limit3_oring_range152w(0) <= below_lower_limit3_oring(1);
	wire_w_exp_and_range8w(0) <= exp_and(0);
	wire_w_exp_and_range14w(0) <= exp_and(1);
	wire_w_exp_and_range19w(0) <= exp_and(2);
	wire_w_exp_and_range24w(0) <= exp_and(3);
	wire_w_exp_and_range29w(0) <= exp_and(4);
	wire_w_exp_and_range34w(0) <= exp_and(5);
	wire_w_exp_and_range39w(0) <= exp_and(6);
	wire_w_exp_bus_range10w(0) <= exp_bus(1);
	wire_w_exp_bus_range15w(0) <= exp_bus(2);
	wire_w_exp_bus_range20w(0) <= exp_bus(3);
	wire_w_exp_bus_range25w(0) <= exp_bus(4);
	wire_w_exp_bus_range30w(0) <= exp_bus(5);
	wire_w_exp_bus_range35w(0) <= exp_bus(6);
	wire_w_exp_bus_range40w(0) <= exp_bus(7);
	wire_w_exp_or_range6w(0) <= exp_or(0);
	wire_w_exp_or_range12w(0) <= exp_or(1);
	wire_w_exp_or_range17w(0) <= exp_or(2);
	wire_w_exp_or_range22w(0) <= exp_or(3);
	wire_w_exp_or_range27w(0) <= exp_or(4);
	wire_w_exp_or_range32w(0) <= exp_or(5);
	wire_w_exp_or_range37w(0) <= exp_or(6);
	wire_w_inv_integer_range250w <= inv_integer(14 DOWNTO 7);
	wire_w_man_bus1_range76w(0) <= man_bus1(0);
	wire_w_man_bus1_range73w(0) <= man_bus1(1);
	wire_w_man_bus1_range70w(0) <= man_bus1(2);
	wire_w_man_bus1_range67w(0) <= man_bus1(3);
	wire_w_man_bus1_range64w(0) <= man_bus1(4);
	wire_w_man_bus1_range61w(0) <= man_bus1(5);
	wire_w_man_bus1_range58w(0) <= man_bus1(6);
	wire_w_man_bus1_range55w(0) <= man_bus1(7);
	wire_w_man_bus1_range52w(0) <= man_bus1(8);
	wire_w_man_bus1_range49w(0) <= man_bus1(9);
	wire_w_man_bus2_range113w(0) <= man_bus2(0);
	wire_w_man_bus2_range83w(0) <= man_bus2(10);
	wire_w_man_bus2_range110w(0) <= man_bus2(1);
	wire_w_man_bus2_range107w(0) <= man_bus2(2);
	wire_w_man_bus2_range104w(0) <= man_bus2(3);
	wire_w_man_bus2_range101w(0) <= man_bus2(4);
	wire_w_man_bus2_range98w(0) <= man_bus2(5);
	wire_w_man_bus2_range95w(0) <= man_bus2(6);
	wire_w_man_bus2_range92w(0) <= man_bus2(7);
	wire_w_man_bus2_range89w(0) <= man_bus2(8);
	wire_w_man_bus2_range86w(0) <= man_bus2(9);
	wire_w_man_or1_range47w(0) <= man_or1(10);
	wire_w_man_or1_range75w(0) <= man_or1(1);
	wire_w_man_or1_range72w(0) <= man_or1(2);
	wire_w_man_or1_range69w(0) <= man_or1(3);
	wire_w_man_or1_range66w(0) <= man_or1(4);
	wire_w_man_or1_range63w(0) <= man_or1(5);
	wire_w_man_or1_range60w(0) <= man_or1(6);
	wire_w_man_or1_range57w(0) <= man_or1(7);
	wire_w_man_or1_range54w(0) <= man_or1(8);
	wire_w_man_or1_range51w(0) <= man_or1(9);
	wire_w_man_or2_range85w(0) <= man_or2(10);
	wire_w_man_or2_range81w(0) <= man_or2(11);
	wire_w_man_or2_range112w(0) <= man_or2(1);
	wire_w_man_or2_range109w(0) <= man_or2(2);
	wire_w_man_or2_range106w(0) <= man_or2(3);
	wire_w_man_or2_range103w(0) <= man_or2(4);
	wire_w_man_or2_range100w(0) <= man_or2(5);
	wire_w_man_or2_range97w(0) <= man_or2(6);
	wire_w_man_or2_range94w(0) <= man_or2(7);
	wire_w_man_or2_range91w(0) <= man_or2(8);
	wire_w_man_or2_range88w(0) <= man_or2(9);
	wire_w_sticky_bus_range200w(0) <= sticky_bus(10);
	wire_w_sticky_bus_range203w(0) <= sticky_bus(11);
	wire_w_sticky_bus_range206w(0) <= sticky_bus(12);
	wire_w_sticky_bus_range209w(0) <= sticky_bus(13);
	wire_w_sticky_bus_range212w(0) <= sticky_bus(14);
	wire_w_sticky_bus_range215w(0) <= sticky_bus(15);
	wire_w_sticky_bus_range218w(0) <= sticky_bus(16);
	wire_w_sticky_bus_range221w(0) <= sticky_bus(17);
	wire_w_sticky_bus_range224w(0) <= sticky_bus(18);
	wire_w_sticky_bus_range227w(0) <= sticky_bus(19);
	wire_w_sticky_bus_range173w(0) <= sticky_bus(1);
	wire_w_sticky_bus_range230w(0) <= sticky_bus(20);
	wire_w_sticky_bus_range233w(0) <= sticky_bus(21);
	wire_w_sticky_bus_range176w(0) <= sticky_bus(2);
	wire_w_sticky_bus_range179w(0) <= sticky_bus(3);
	wire_w_sticky_bus_range182w(0) <= sticky_bus(4);
	wire_w_sticky_bus_range185w(0) <= sticky_bus(5);
	wire_w_sticky_bus_range188w(0) <= sticky_bus(6);
	wire_w_sticky_bus_range191w(0) <= sticky_bus(7);
	wire_w_sticky_bus_range194w(0) <= sticky_bus(8);
	wire_w_sticky_bus_range197w(0) <= sticky_bus(9);
	wire_w_sticky_or_range171w(0) <= sticky_or(0);
	wire_w_sticky_or_range202w(0) <= sticky_or(10);
	wire_w_sticky_or_range205w(0) <= sticky_or(11);
	wire_w_sticky_or_range208w(0) <= sticky_or(12);
	wire_w_sticky_or_range211w(0) <= sticky_or(13);
	wire_w_sticky_or_range214w(0) <= sticky_or(14);
	wire_w_sticky_or_range217w(0) <= sticky_or(15);
	wire_w_sticky_or_range220w(0) <= sticky_or(16);
	wire_w_sticky_or_range223w(0) <= sticky_or(17);
	wire_w_sticky_or_range226w(0) <= sticky_or(18);
	wire_w_sticky_or_range229w(0) <= sticky_or(19);
	wire_w_sticky_or_range175w(0) <= sticky_or(1);
	wire_w_sticky_or_range232w(0) <= sticky_or(20);
	wire_w_sticky_or_range178w(0) <= sticky_or(2);
	wire_w_sticky_or_range181w(0) <= sticky_or(3);
	wire_w_sticky_or_range184w(0) <= sticky_or(4);
	wire_w_sticky_or_range187w(0) <= sticky_or(5);
	wire_w_sticky_or_range190w(0) <= sticky_or(6);
	wire_w_sticky_or_range193w(0) <= sticky_or(7);
	wire_w_sticky_or_range196w(0) <= sticky_or(8);
	wire_w_sticky_or_range199w(0) <= sticky_or(9);
	wire_altbarrel_shift2_distance <= wire_w_lg_w_lg_barrel_direction_negative164w165w;
	loop44 : FOR i IN 0 TO 5 GENERATE 
		wire_w_lg_w_lg_barrel_direction_negative164w165w(i) <= wire_w_lg_barrel_direction_negative164w(i) OR wire_w_lg_w_lg_barrel_direction_negative162w163w(i);
	END GENERATE loop44;
	altbarrel_shift2 :  fp32_signed16_conv_altbarrel_shift_i4h
	  PORT MAP ( 
		aclr => aclr,
		clk_en => clk_en,
		clock => clock,
		data => barrel_mantissa_input,
		direction => barrel_direction_negative,
		distance => wire_altbarrel_shift2_distance,
		result => wire_altbarrel_shift2_result
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN added_power2_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN added_power2_reg <= wire_add_sub1_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_direction_negative_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_direction_negative_reg <= wire_power2_value_w_result_range146w(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit2_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit2_reg1 <= below_lower_limit2_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit2_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit2_reg2 <= below_lower_limit2_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit2_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit2_reg3 <= below_lower_limit2_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit2_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit2_reg4 <= below_lower_limit2_reg3;
			END IF;
		END IF;
	END PROCESS;
	wire_below_lower_limit2_reg4_w_lg_q288w(0) <= below_lower_limit2_reg4 AND wire_border_lower_limit_reg4_w_lg_q287w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit3_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit3_reg1 <= below_lower_limit3_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit3_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit3_reg2 <= below_lower_limit3_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit3_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit3_reg3 <= below_lower_limit3_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit3_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit3_reg4 <= below_lower_limit3_reg3;
			END IF;
		END IF;
	END PROCESS;
	wire_below_lower_limit3_reg4_w_lg_q292w(0) <= below_lower_limit3_reg4 AND wire_w_lg_zero_input_w291w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN border_lower_limit_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN border_lower_limit_reg1 <= wire_below_lower_limit2_aeb;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN border_lower_limit_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN border_lower_limit_reg2 <= border_lower_limit_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN border_lower_limit_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN border_lower_limit_reg3 <= border_lower_limit_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN border_lower_limit_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN border_lower_limit_reg4 <= border_lower_limit_reg3;
			END IF;
		END IF;
	END PROCESS;
	wire_border_lower_limit_reg4_w_lg_q287w(0) <= NOT border_lower_limit_reg4;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dataa_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dataa_reg <= dataa;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN equal_upper_limit_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN equal_upper_limit_reg1 <= equal_upper_limit_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN equal_upper_limit_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN equal_upper_limit_reg2 <= equal_upper_limit_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN equal_upper_limit_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN equal_upper_limit_reg3 <= equal_upper_limit_reg2;
			END IF;
		END IF;
	END PROCESS;
	wire_equal_upper_limit_reg3_w_lg_q252w(0) <= equal_upper_limit_reg3 AND wire_int_or_reg3_w_lg_q251w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exceed_upper_limit_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exceed_upper_limit_reg1 <= exceed_upper_limit_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exceed_upper_limit_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exceed_upper_limit_reg2 <= exceed_upper_limit_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exceed_upper_limit_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exceed_upper_limit_reg3 <= exceed_upper_limit_reg2;
			END IF;
		END IF;
	END PROCESS;
	wire_exceed_upper_limit_reg3_w_lg_q253w(0) <= exceed_upper_limit_reg3 OR wire_equal_upper_limit_reg3_w_lg_q252w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exceed_upper_limit_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exceed_upper_limit_reg4 <= upper_limit_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_and_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_and_reg1 <= exp_and_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_and_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_and_reg2 <= exp_and_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_and_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_and_reg3 <= exp_and_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_and_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_and_reg4 <= exp_and_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_or_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_or_reg1 <= exp_or_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_or_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_or_reg2 <= exp_or_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_or_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_or_reg3 <= exp_or_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_or_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_or_reg4 <= exp_or_reg3;
			END IF;
		END IF;
	END PROCESS;
	wire_exp_or_reg4_w_lg_q118w(0) <= NOT exp_or_reg4;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN int_or1_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN int_or1_reg1 <= int_or1_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN int_or2_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN int_or2_reg1 <= int_or2_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN int_or_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN int_or_reg2 <= (int_or1_reg1 OR int_or2_reg1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN int_or_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN int_or_reg3 <= int_or_reg2;
			END IF;
		END IF;
	END PROCESS;
	wire_int_or_reg3_w_lg_q251w(0) <= int_or_reg3 OR add_1_w;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN integer_result_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN integer_result_reg <= integer_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN integer_rounded_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN integer_rounded_reg <= integer_rounded;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lowest_int_sel_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lowest_int_sel_reg <= lowest_integer_selector;
			END IF;
		END IF;
	END PROCESS;
	wire_lowest_int_sel_reg_w_lg_q289w(0) <= NOT lowest_int_sel_reg;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_or1_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_or1_reg1 <= man_or1_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_or2_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_or2_reg1 <= man_or2_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_or_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_or_reg2 <= man_or_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_or_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_or_reg3 <= man_or_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_or_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_or_reg4 <= man_or_reg3;
			END IF;
		END IF;
	END PROCESS;
	wire_man_or_reg4_w_lg_q120w(0) <= NOT man_or_reg4;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mantissa_input_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mantissa_input_reg <= mantissa_input;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN max_shift_exceeder_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN max_shift_exceeder_reg <= more_than_max_shift_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN max_shift_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN max_shift_reg <= wire_max_shift_compare_agb;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_reg <= nan_input_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN overflow_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN overflow_reg <= exceed_limit_exceeders;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN power2_value_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN power2_value_reg <= power2_value_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_input_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_input_reg1 <= sign_input;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_input_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_input_reg2 <= sign_input_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_input_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_input_reg3 <= sign_input_reg2;
			END IF;
		END IF;
	END PROCESS;
	wire_sign_input_reg3_w_lg_q254w(0) <= sign_input_reg3 AND wire_exceed_upper_limit_reg3_w_lg_q253w(0);
	wire_sign_input_reg3_w_lg_q256w(0) <= NOT sign_input_reg3;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_input_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_input_reg4 <= sign_input_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN underflow_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN underflow_reg <= lower_limit_selector;
			END IF;
		END IF;
	END PROCESS;
	wire_add_1_adder_datab <= "000000000000001";
	add_1_adder :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 15,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		cout => wire_add_1_adder_cout,
		dataa => integer_pre_round,
		datab => wire_add_1_adder_datab,
		result => wire_add_1_adder_result
	  );
	wire_add_sub1_datab <= "000001";
	add_sub1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 6,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => power2_value_reg,
		datab => wire_add_sub1_datab,
		result => wire_add_sub1_result
	  );
	loop45 : FOR i IN 0 TO 7 GENERATE 
		wire_add_sub3_w_lg_w_lg_cout263w264w(i) <= wire_add_sub3_w_lg_cout263w(0) AND wire_w_inv_integer_range250w(i);
	END GENERATE loop45;
	loop46 : FOR i IN 0 TO 7 GENERATE 
		wire_add_sub3_w_lg_cout262w(i) <= wire_add_sub3_cout AND wire_add_sub4_result(i);
	END GENERATE loop46;
	wire_add_sub3_w_lg_cout263w(0) <= NOT wire_add_sub3_cout;
	wire_add_sub3_datab <= "0000001";
	add_sub3 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 7,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		cout => wire_add_sub3_cout,
		dataa => inv_integer(6 DOWNTO 0),
		datab => wire_add_sub3_datab,
		result => wire_add_sub3_result
	  );
	wire_add_sub4_datab <= "00000001";
	add_sub4 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 8,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => inv_integer(14 DOWNTO 7),
		datab => wire_add_sub4_datab,
		result => wire_add_sub4_result
	  );
	wire_barrel_direction_invert_dataa <= (OTHERS => '0');
	barrel_direction_invert :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_WIDTH => 6,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => wire_barrel_direction_invert_dataa,
		datab => power2_value_reg,
		result => wire_barrel_direction_invert_result
	  );
	wire_power2_value_w_lg_w_result_range146w154w(0) <= wire_power2_value_w_result_range146w(0) AND wire_w_below_lower_limit3_oring_range152w(0);
	wire_power2_value_w_lg_w_lg_w_result_range146w154w155w(0) <= wire_power2_value_w_lg_w_result_range146w154w(0) OR power2_value_overflow_w;
	wire_power2_value_w_result_range128w(0) <= wire_power2_value_result(1);
	wire_power2_value_w_result_range131w(0) <= wire_power2_value_result(2);
	wire_power2_value_w_result_range134w(0) <= wire_power2_value_result(3);
	wire_power2_value_w_result_range137w(0) <= wire_power2_value_result(4);
	wire_power2_value_w_result_range140w(0) <= wire_power2_value_result(5);
	wire_power2_value_w_result_range143w(0) <= wire_power2_value_result(6);
	wire_power2_value_w_result_range146w(0) <= wire_power2_value_result(7);
	power2_value :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => exponent_input,
		datab => shift_value_w,
		overflow => wire_power2_value_overflow,
		result => wire_power2_value_result
	  );
	below_lower_limit1 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		aeb => wire_below_lower_limit1_aeb,
		dataa => exponent_input,
		datab => bias_value_less_1_w
	  );
	below_lower_limit2 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		aeb => wire_below_lower_limit2_aeb,
		alb => wire_below_lower_limit2_alb,
		dataa => exponent_input,
		datab => shift_value_w
	  );
	exceed_upper_limit :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		aeb => wire_exceed_upper_limit_aeb,
		agb => wire_exceed_upper_limit_agb,
		dataa => padded_exponent_input,
		datab => const_bias_value_add_width_res_w
	  );
	max_shift_compare :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		agb => wire_max_shift_compare_agb,
		dataa => added_power2_reg,
		datab => max_shift_w
	  );

 END RTL; --fp32_signed16_conv_altfp_convert_46p
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY fp32_signed16_conv IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		dataa		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		nan		: OUT STD_LOGIC ;
		overflow		: OUT STD_LOGIC ;
		result		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		underflow		: OUT STD_LOGIC 
	);
END fp32_signed16_conv;


ARCHITECTURE RTL OF fp32_signed16_conv IS

	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC ;
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC ;



	COMPONENT fp32_signed16_conv_altfp_convert_46p
	PORT (
			clock	: IN STD_LOGIC ;
			dataa	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			nan	: OUT STD_LOGIC ;
			overflow	: OUT STD_LOGIC ;
			result	: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
			underflow	: OUT STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	nan    <= sub_wire0;
	overflow    <= sub_wire1;
	result    <= sub_wire2(15 DOWNTO 0);
	underflow    <= sub_wire3;

	fp32_signed16_conv_altfp_convert_46p_component : fp32_signed16_conv_altfp_convert_46p
	PORT MAP (
		clock => clock,
		dataa => dataa,
		nan => sub_wire0,
		overflow => sub_wire1,
		result => sub_wire2,
		underflow => sub_wire3
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altfp_convert"
-- Retrieval info: CONSTANT: OPERATION STRING "FLOAT2FIXED"
-- Retrieval info: CONSTANT: ROUNDING STRING "TO_NEAREST"
-- Retrieval info: CONSTANT: WIDTH_DATA NUMERIC "32"
-- Retrieval info: CONSTANT: WIDTH_EXP_INPUT NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_EXP_OUTPUT NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_INT NUMERIC "4"
-- Retrieval info: CONSTANT: WIDTH_MAN_INPUT NUMERIC "23"
-- Retrieval info: CONSTANT: WIDTH_MAN_OUTPUT NUMERIC "23"
-- Retrieval info: CONSTANT: WIDTH_RESULT NUMERIC "16"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: USED_PORT: dataa 0 0 32 0 INPUT NODEFVAL "dataa[31..0]"
-- Retrieval info: CONNECT: @dataa 0 0 32 0 dataa 0 0 32 0
-- Retrieval info: USED_PORT: nan 0 0 0 0 OUTPUT NODEFVAL "nan"
-- Retrieval info: CONNECT: nan 0 0 0 0 @nan 0 0 0 0
-- Retrieval info: USED_PORT: overflow 0 0 0 0 OUTPUT NODEFVAL "overflow"
-- Retrieval info: CONNECT: overflow 0 0 0 0 @overflow 0 0 0 0
-- Retrieval info: USED_PORT: result 0 0 16 0 OUTPUT NODEFVAL "result[15..0]"
-- Retrieval info: CONNECT: result 0 0 16 0 @result 0 0 16 0
-- Retrieval info: USED_PORT: underflow 0 0 0 0 OUTPUT NODEFVAL "underflow"
-- Retrieval info: CONNECT: underflow 0 0 0 0 @underflow 0 0 0 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL fp32_signed16_conv.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fp32_signed16_conv.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fp32_signed16_conv.bsf TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fp32_signed16_conv_inst.vhd TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fp32_signed16_conv.inc TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fp32_signed16_conv.cmp TRUE TRUE
-- Retrieval info: LIB_FILE: lpm
