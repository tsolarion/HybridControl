LVDS_ALT_inst : LVDS_ALT PORT MAP (
		tx_in	 => tx_in_sig,
		tx_inclock	 => tx_inclock_sig,
		tx_syncclock	 => tx_syncclock_sig,
		tx_out	 => tx_out_sig
	);
